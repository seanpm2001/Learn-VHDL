-- this is a single line VHDL comment
/*
    this is a block comment (in VHDL-2008 and later)
*/
